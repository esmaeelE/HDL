module ANDGate (output wire Y, input wire A, input wire B);
            assign Y = A & B;
endmodule
        