// hello module definition in verilog

module hello;
  initial
    begin
      $display("Hello, World");
      $finish ;
    end
endmodule



